// qsys_system.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module qsys_system (
		input  wire        clk_clk,             //          clk.clk
		output wire [7:0]  control_bits_export, // control_bits.export
		output wire [7:0]  dac_div_export,      //      dac_div.export
		output wire [7:0]  dac_gain_export,     //     dac_gain.export
		output wire [5:0]  gain_ctrl_export,    //    gain_ctrl.export
		input  wire [15:0] lia_1_x_export,      //      lia_1_x.export
		input  wire [15:0] lia_1_y_export,      //      lia_1_y.export
		output wire [19:0] phase_incr_1_export, // phase_incr_1.export
		output wire [19:0] phase_incr_2_export, // phase_incr_2.export
		output wire [19:0] phase_incr_3_export, // phase_incr_3.export
		output wire [19:0] phase_incr_4_export, // phase_incr_4.export
		output wire [19:0] phase_incr_5_export, // phase_incr_5.export
		output wire [19:0] phase_incr_6_export, // phase_incr_6.export
		output wire [19:0] phase_incr_7_export, // phase_incr_7.export
		output wire [19:0] phase_incr_8_export, // phase_incr_8.export
		output wire [19:0] phase_offs_1_export, // phase_offs_1.export
		output wire [19:0] phase_offs_2_export, // phase_offs_2.export
		output wire [19:0] phase_offs_3_export, // phase_offs_3.export
		output wire [19:0] phase_offs_4_export, // phase_offs_4.export
		output wire [19:0] phase_offs_5_export, // phase_offs_5.export
		output wire [19:0] phase_offs_6_export, // phase_offs_6.export
		output wire [19:0] phase_offs_7_export, // phase_offs_7.export
		output wire [19:0] phase_offs_8_export, // phase_offs_8.export
		input  wire        reset_reset_n,       //        reset.reset_n
		output wire        resetrequest_reset   // resetrequest.reset
	);

	wire  [31:0] bfm_master_m0_readdata;                             // mm_interconnect_0:bfm_master_m0_readdata -> bfm_master:avm_readdata
	wire         bfm_master_m0_waitrequest;                          // mm_interconnect_0:bfm_master_m0_waitrequest -> bfm_master:avm_waitrequest
	wire  [31:0] bfm_master_m0_address;                              // bfm_master:avm_address -> mm_interconnect_0:bfm_master_m0_address
	wire         bfm_master_m0_read;                                 // bfm_master:avm_read -> mm_interconnect_0:bfm_master_m0_read
	wire   [3:0] bfm_master_m0_byteenable;                           // bfm_master:avm_byteenable -> mm_interconnect_0:bfm_master_m0_byteenable
	wire         bfm_master_m0_readdatavalid;                        // mm_interconnect_0:bfm_master_m0_readdatavalid -> bfm_master:avm_readdatavalid
	wire  [31:0] bfm_master_m0_writedata;                            // bfm_master:avm_writedata -> mm_interconnect_0:bfm_master_m0_writedata
	wire         bfm_master_m0_write;                                // bfm_master:avm_write -> mm_interconnect_0:bfm_master_m0_write
	wire  [31:0] jtag_master_master_readdata;                        // mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	wire         jtag_master_master_waitrequest;                     // mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	wire  [31:0] jtag_master_master_address;                         // jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	wire         jtag_master_master_read;                            // jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	wire   [3:0] jtag_master_master_byteenable;                      // jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	wire         jtag_master_master_readdatavalid;                   // mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	wire         jtag_master_master_write;                           // jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	wire  [31:0] jtag_master_master_writedata;                       // jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	wire         mm_interconnect_0_nco_freq_control_1_s1_chipselect; // mm_interconnect_0:nco_freq_control_1_s1_chipselect -> nco_freq_control_1:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_control_1_s1_readdata;   // nco_freq_control_1:readdata -> mm_interconnect_0:nco_freq_control_1_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_control_1_s1_address;    // mm_interconnect_0:nco_freq_control_1_s1_address -> nco_freq_control_1:address
	wire         mm_interconnect_0_nco_freq_control_1_s1_write;      // mm_interconnect_0:nco_freq_control_1_s1_write -> nco_freq_control_1:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_control_1_s1_writedata;  // mm_interconnect_0:nco_freq_control_1_s1_writedata -> nco_freq_control_1:writedata
	wire         mm_interconnect_0_nco_freq_control_2_s1_chipselect; // mm_interconnect_0:nco_freq_control_2_s1_chipselect -> nco_freq_control_2:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_control_2_s1_readdata;   // nco_freq_control_2:readdata -> mm_interconnect_0:nco_freq_control_2_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_control_2_s1_address;    // mm_interconnect_0:nco_freq_control_2_s1_address -> nco_freq_control_2:address
	wire         mm_interconnect_0_nco_freq_control_2_s1_write;      // mm_interconnect_0:nco_freq_control_2_s1_write -> nco_freq_control_2:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_control_2_s1_writedata;  // mm_interconnect_0:nco_freq_control_2_s1_writedata -> nco_freq_control_2:writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;         // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;           // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_ram_s1_address;            // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;         // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;              // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;          // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;              // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_1_s1_chipselect -> nco_phase_ctrl_1:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_1_s1_readdata;     // nco_phase_ctrl_1:readdata -> mm_interconnect_0:nco_phase_ctrl_1_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_1_s1_address;      // mm_interconnect_0:nco_phase_ctrl_1_s1_address -> nco_phase_ctrl_1:address
	wire         mm_interconnect_0_nco_phase_ctrl_1_s1_write;        // mm_interconnect_0:nco_phase_ctrl_1_s1_write -> nco_phase_ctrl_1:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_1_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_1_s1_writedata -> nco_phase_ctrl_1:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_2_s1_chipselect -> nco_phase_ctrl_2:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_2_s1_readdata;     // nco_phase_ctrl_2:readdata -> mm_interconnect_0:nco_phase_ctrl_2_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_2_s1_address;      // mm_interconnect_0:nco_phase_ctrl_2_s1_address -> nco_phase_ctrl_2:address
	wire         mm_interconnect_0_nco_phase_ctrl_2_s1_write;        // mm_interconnect_0:nco_phase_ctrl_2_s1_write -> nco_phase_ctrl_2:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_2_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_2_s1_writedata -> nco_phase_ctrl_2:writedata
	wire         mm_interconnect_0_gain_controller_s1_chipselect;    // mm_interconnect_0:gain_controller_s1_chipselect -> gain_controller:chipselect
	wire  [31:0] mm_interconnect_0_gain_controller_s1_readdata;      // gain_controller:readdata -> mm_interconnect_0:gain_controller_s1_readdata
	wire   [1:0] mm_interconnect_0_gain_controller_s1_address;       // mm_interconnect_0:gain_controller_s1_address -> gain_controller:address
	wire         mm_interconnect_0_gain_controller_s1_write;         // mm_interconnect_0:gain_controller_s1_write -> gain_controller:write_n
	wire  [31:0] mm_interconnect_0_gain_controller_s1_writedata;     // mm_interconnect_0:gain_controller_s1_writedata -> gain_controller:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_3_s1_chipselect -> nco_freq_ctrl_3:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_3_s1_readdata;      // nco_freq_ctrl_3:readdata -> mm_interconnect_0:nco_freq_ctrl_3_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_3_s1_address;       // mm_interconnect_0:nco_freq_ctrl_3_s1_address -> nco_freq_ctrl_3:address
	wire         mm_interconnect_0_nco_freq_ctrl_3_s1_write;         // mm_interconnect_0:nco_freq_ctrl_3_s1_write -> nco_freq_ctrl_3:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_3_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_3_s1_writedata -> nco_freq_ctrl_3:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_4_s1_chipselect -> nco_freq_ctrl_4:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_4_s1_readdata;      // nco_freq_ctrl_4:readdata -> mm_interconnect_0:nco_freq_ctrl_4_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_4_s1_address;       // mm_interconnect_0:nco_freq_ctrl_4_s1_address -> nco_freq_ctrl_4:address
	wire         mm_interconnect_0_nco_freq_ctrl_4_s1_write;         // mm_interconnect_0:nco_freq_ctrl_4_s1_write -> nco_freq_ctrl_4:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_4_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_4_s1_writedata -> nco_freq_ctrl_4:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_5_s1_chipselect -> nco_freq_ctrl_5:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_5_s1_readdata;      // nco_freq_ctrl_5:readdata -> mm_interconnect_0:nco_freq_ctrl_5_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_5_s1_address;       // mm_interconnect_0:nco_freq_ctrl_5_s1_address -> nco_freq_ctrl_5:address
	wire         mm_interconnect_0_nco_freq_ctrl_5_s1_write;         // mm_interconnect_0:nco_freq_ctrl_5_s1_write -> nco_freq_ctrl_5:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_5_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_5_s1_writedata -> nco_freq_ctrl_5:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_6_s1_chipselect -> nco_freq_ctrl_6:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_6_s1_readdata;      // nco_freq_ctrl_6:readdata -> mm_interconnect_0:nco_freq_ctrl_6_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_6_s1_address;       // mm_interconnect_0:nco_freq_ctrl_6_s1_address -> nco_freq_ctrl_6:address
	wire         mm_interconnect_0_nco_freq_ctrl_6_s1_write;         // mm_interconnect_0:nco_freq_ctrl_6_s1_write -> nco_freq_ctrl_6:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_6_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_6_s1_writedata -> nco_freq_ctrl_6:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_7_s1_chipselect -> nco_freq_ctrl_7:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_7_s1_readdata;      // nco_freq_ctrl_7:readdata -> mm_interconnect_0:nco_freq_ctrl_7_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_7_s1_address;       // mm_interconnect_0:nco_freq_ctrl_7_s1_address -> nco_freq_ctrl_7:address
	wire         mm_interconnect_0_nco_freq_ctrl_7_s1_write;         // mm_interconnect_0:nco_freq_ctrl_7_s1_write -> nco_freq_ctrl_7:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_7_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_7_s1_writedata -> nco_freq_ctrl_7:writedata
	wire         mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect;    // mm_interconnect_0:nco_freq_ctrl_8_s1_chipselect -> nco_freq_ctrl_8:chipselect
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_8_s1_readdata;      // nco_freq_ctrl_8:readdata -> mm_interconnect_0:nco_freq_ctrl_8_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_freq_ctrl_8_s1_address;       // mm_interconnect_0:nco_freq_ctrl_8_s1_address -> nco_freq_ctrl_8:address
	wire         mm_interconnect_0_nco_freq_ctrl_8_s1_write;         // mm_interconnect_0:nco_freq_ctrl_8_s1_write -> nco_freq_ctrl_8:write_n
	wire  [31:0] mm_interconnect_0_nco_freq_ctrl_8_s1_writedata;     // mm_interconnect_0:nco_freq_ctrl_8_s1_writedata -> nco_freq_ctrl_8:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_3_s1_chipselect -> nco_phase_ctrl_3:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_3_s1_readdata;     // nco_phase_ctrl_3:readdata -> mm_interconnect_0:nco_phase_ctrl_3_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_3_s1_address;      // mm_interconnect_0:nco_phase_ctrl_3_s1_address -> nco_phase_ctrl_3:address
	wire         mm_interconnect_0_nco_phase_ctrl_3_s1_write;        // mm_interconnect_0:nco_phase_ctrl_3_s1_write -> nco_phase_ctrl_3:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_3_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_3_s1_writedata -> nco_phase_ctrl_3:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_4_s1_chipselect -> nco_phase_ctrl_4:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_4_s1_readdata;     // nco_phase_ctrl_4:readdata -> mm_interconnect_0:nco_phase_ctrl_4_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_4_s1_address;      // mm_interconnect_0:nco_phase_ctrl_4_s1_address -> nco_phase_ctrl_4:address
	wire         mm_interconnect_0_nco_phase_ctrl_4_s1_write;        // mm_interconnect_0:nco_phase_ctrl_4_s1_write -> nco_phase_ctrl_4:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_4_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_4_s1_writedata -> nco_phase_ctrl_4:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_5_s1_chipselect -> nco_phase_ctrl_5:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_5_s1_readdata;     // nco_phase_ctrl_5:readdata -> mm_interconnect_0:nco_phase_ctrl_5_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_5_s1_address;      // mm_interconnect_0:nco_phase_ctrl_5_s1_address -> nco_phase_ctrl_5:address
	wire         mm_interconnect_0_nco_phase_ctrl_5_s1_write;        // mm_interconnect_0:nco_phase_ctrl_5_s1_write -> nco_phase_ctrl_5:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_5_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_5_s1_writedata -> nco_phase_ctrl_5:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_6_s1_chipselect -> nco_phase_ctrl_6:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_6_s1_readdata;     // nco_phase_ctrl_6:readdata -> mm_interconnect_0:nco_phase_ctrl_6_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_6_s1_address;      // mm_interconnect_0:nco_phase_ctrl_6_s1_address -> nco_phase_ctrl_6:address
	wire         mm_interconnect_0_nco_phase_ctrl_6_s1_write;        // mm_interconnect_0:nco_phase_ctrl_6_s1_write -> nco_phase_ctrl_6:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_6_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_6_s1_writedata -> nco_phase_ctrl_6:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_7_s1_chipselect -> nco_phase_ctrl_7:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_7_s1_readdata;     // nco_phase_ctrl_7:readdata -> mm_interconnect_0:nco_phase_ctrl_7_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_7_s1_address;      // mm_interconnect_0:nco_phase_ctrl_7_s1_address -> nco_phase_ctrl_7:address
	wire         mm_interconnect_0_nco_phase_ctrl_7_s1_write;        // mm_interconnect_0:nco_phase_ctrl_7_s1_write -> nco_phase_ctrl_7:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_7_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_7_s1_writedata -> nco_phase_ctrl_7:writedata
	wire         mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect;   // mm_interconnect_0:nco_phase_ctrl_8_s1_chipselect -> nco_phase_ctrl_8:chipselect
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_8_s1_readdata;     // nco_phase_ctrl_8:readdata -> mm_interconnect_0:nco_phase_ctrl_8_s1_readdata
	wire   [1:0] mm_interconnect_0_nco_phase_ctrl_8_s1_address;      // mm_interconnect_0:nco_phase_ctrl_8_s1_address -> nco_phase_ctrl_8:address
	wire         mm_interconnect_0_nco_phase_ctrl_8_s1_write;        // mm_interconnect_0:nco_phase_ctrl_8_s1_write -> nco_phase_ctrl_8:write_n
	wire  [31:0] mm_interconnect_0_nco_phase_ctrl_8_s1_writedata;    // mm_interconnect_0:nco_phase_ctrl_8_s1_writedata -> nco_phase_ctrl_8:writedata
	wire  [31:0] mm_interconnect_0_lia_1_x_s1_readdata;              // lia_1_x:readdata -> mm_interconnect_0:lia_1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_lia_1_x_s1_address;               // mm_interconnect_0:lia_1_x_s1_address -> lia_1_x:address
	wire  [31:0] mm_interconnect_0_lia_1_y_s1_readdata;              // lia_1_y:readdata -> mm_interconnect_0:lia_1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_lia_1_y_s1_address;               // mm_interconnect_0:lia_1_y_s1_address -> lia_1_y:address
	wire         mm_interconnect_0_dac_gain_s1_chipselect;           // mm_interconnect_0:dac_gain_s1_chipselect -> dac_gain:chipselect
	wire  [31:0] mm_interconnect_0_dac_gain_s1_readdata;             // dac_gain:readdata -> mm_interconnect_0:dac_gain_s1_readdata
	wire   [1:0] mm_interconnect_0_dac_gain_s1_address;              // mm_interconnect_0:dac_gain_s1_address -> dac_gain:address
	wire         mm_interconnect_0_dac_gain_s1_write;                // mm_interconnect_0:dac_gain_s1_write -> dac_gain:write_n
	wire  [31:0] mm_interconnect_0_dac_gain_s1_writedata;            // mm_interconnect_0:dac_gain_s1_writedata -> dac_gain:writedata
	wire         mm_interconnect_0_dac_div_s1_chipselect;            // mm_interconnect_0:dac_div_s1_chipselect -> dac_div:chipselect
	wire  [31:0] mm_interconnect_0_dac_div_s1_readdata;              // dac_div:readdata -> mm_interconnect_0:dac_div_s1_readdata
	wire   [1:0] mm_interconnect_0_dac_div_s1_address;               // mm_interconnect_0:dac_div_s1_address -> dac_div:address
	wire         mm_interconnect_0_dac_div_s1_write;                 // mm_interconnect_0:dac_div_s1_write -> dac_div:write_n
	wire  [31:0] mm_interconnect_0_dac_div_s1_writedata;             // mm_interconnect_0:dac_div_s1_writedata -> dac_div:writedata
	wire         mm_interconnect_0_control_bits_s1_chipselect;       // mm_interconnect_0:control_bits_s1_chipselect -> control_bits:chipselect
	wire  [31:0] mm_interconnect_0_control_bits_s1_readdata;         // control_bits:readdata -> mm_interconnect_0:control_bits_s1_readdata
	wire   [1:0] mm_interconnect_0_control_bits_s1_address;          // mm_interconnect_0:control_bits_s1_address -> control_bits:address
	wire         mm_interconnect_0_control_bits_s1_write;            // mm_interconnect_0:control_bits_s1_write -> control_bits:write_n
	wire  [31:0] mm_interconnect_0_control_bits_s1_writedata;        // mm_interconnect_0:control_bits_s1_writedata -> control_bits:writedata
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [bfm_master:reset, control_bits:reset_n, dac_div:reset_n, dac_gain:reset_n, gain_controller:reset_n, lia_1_x:reset_n, lia_1_y:reset_n, mm_interconnect_0:bfm_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, nco_freq_control_1:reset_n, nco_freq_control_2:reset_n, nco_freq_ctrl_3:reset_n, nco_freq_ctrl_4:reset_n, nco_freq_ctrl_5:reset_n, nco_freq_ctrl_6:reset_n, nco_freq_ctrl_7:reset_n, nco_freq_ctrl_8:reset_n, nco_phase_ctrl_1:reset_n, nco_phase_ctrl_2:reset_n, nco_phase_ctrl_3:reset_n, nco_phase_ctrl_4:reset_n, nco_phase_ctrl_5:reset_n, nco_phase_ctrl_6:reset_n, nco_phase_ctrl_7:reset_n, nco_phase_ctrl_8:reset_n, onchip_ram:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [onchip_ram:reset_req, rst_translator:reset_req_in]

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (32),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (4),
		.AV_BURSTCOUNT_W            (3),
		.AV_READRESPONSE_W          (8),
		.AV_WRITERESPONSE_W         (8),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (1),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (1),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (1),
		.AV_MAX_PENDING_READS       (0),
		.AV_MAX_PENDING_WRITES      (0),
		.AV_FIX_READ_LATENCY        (1),
		.AV_READ_WAIT_TIME          (1),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0),
		.VHDL_ID                    (0)
	) bfm_master (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.avm_address            (bfm_master_m0_address),          //        m0.address
		.avm_readdata           (bfm_master_m0_readdata),         //          .readdata
		.avm_writedata          (bfm_master_m0_writedata),        //          .writedata
		.avm_waitrequest        (bfm_master_m0_waitrequest),      //          .waitrequest
		.avm_write              (bfm_master_m0_write),            //          .write
		.avm_read               (bfm_master_m0_read),             //          .read
		.avm_byteenable         (bfm_master_m0_byteenable),       //          .byteenable
		.avm_readdatavalid      (bfm_master_m0_readdatavalid),    //          .readdatavalid
		.avm_burstcount         (),                               // (terminated)
		.avm_begintransfer      (),                               // (terminated)
		.avm_beginbursttransfer (),                               // (terminated)
		.avm_arbiterlock        (),                               // (terminated)
		.avm_lock               (),                               // (terminated)
		.avm_debugaccess        (),                               // (terminated)
		.avm_transactionid      (),                               // (terminated)
		.avm_readid             (8'b00000000),                    // (terminated)
		.avm_writeid            (8'b00000000),                    // (terminated)
		.avm_clken              (),                               // (terminated)
		.avm_response           (2'b00),                          // (terminated)
		.avm_writeresponsevalid (1'b0),                           // (terminated)
		.avm_readresponse       (8'b00000000),                    // (terminated)
		.avm_writeresponse      (8'b00000000)                     // (terminated)
	);

	qsys_system_control_bits control_bits (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_control_bits_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_control_bits_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_control_bits_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_control_bits_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_control_bits_s1_readdata),   //                    .readdata
		.out_port   (control_bits_export)                           // external_connection.export
	);

	qsys_system_control_bits dac_div (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_dac_div_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dac_div_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dac_div_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dac_div_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dac_div_s1_readdata),   //                    .readdata
		.out_port   (dac_div_export)                           // external_connection.export
	);

	qsys_system_dac_gain dac_gain (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_dac_gain_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dac_gain_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dac_gain_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dac_gain_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dac_gain_s1_readdata),   //                    .readdata
		.out_port   (dac_gain_export)                           // external_connection.export
	);

	qsys_system_gain_controller gain_controller (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_gain_controller_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gain_controller_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gain_controller_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gain_controller_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gain_controller_s1_readdata),   //                    .readdata
		.out_port   (gain_ctrl_export)                                 // external_connection.export
	);

	qsys_system_jtag_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (clk_clk),                          //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                   //    clk_reset.reset
		.master_address       (jtag_master_master_address),       //       master.address
		.master_readdata      (jtag_master_master_readdata),      //             .readdata
		.master_read          (jtag_master_master_read),          //             .read
		.master_write         (jtag_master_master_write),         //             .write
		.master_writedata     (jtag_master_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),    //             .byteenable
		.master_reset_reset   (resetrequest_reset)                // master_reset.reset
	);

	qsys_system_lia_1_x lia_1_x (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_lia_1_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lia_1_x_s1_readdata), //                    .readdata
		.in_port  (lia_1_x_export)                         // external_connection.export
	);

	qsys_system_lia_1_x lia_1_y (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_lia_1_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_lia_1_y_s1_readdata), //                    .readdata
		.in_port  (lia_1_y_export)                         // external_connection.export
	);

	qsys_system_nco_freq_control_1 nco_freq_control_1 (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_control_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_control_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_control_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_control_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_control_1_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_1_export)                                 // external_connection.export
	);

	qsys_system_nco_freq_control_1 nco_freq_control_2 (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_control_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_control_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_control_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_control_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_control_2_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_2_export)                                 // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_3 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_3_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_3_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_4 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_4_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_4_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_5 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_5_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_5_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_6 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_6_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_6_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_7 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_7_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_7_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_freq_ctrl_8 (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_nco_freq_ctrl_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_freq_ctrl_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_freq_ctrl_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_freq_ctrl_8_s1_readdata),   //                    .readdata
		.out_port   (phase_incr_8_export)                              // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_1 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_1_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_1_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_2 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_2_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_2_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_3 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_3_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_3_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_4 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_4_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_4_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_5 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_5_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_5_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_6 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_6_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_6_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_7 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_7_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_7_export)                               // external_connection.export
	);

	qsys_system_nco_freq_ctrl_3 nco_phase_ctrl_8 (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_nco_phase_ctrl_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_nco_phase_ctrl_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_nco_phase_ctrl_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_nco_phase_ctrl_8_s1_readdata),   //                    .readdata
		.out_port   (phase_offs_8_export)                               // external_connection.export
	);

	qsys_system_onchip_ram onchip_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	qsys_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                       (clk_clk),                                            //                                     clk_clk.clk
		.bfm_master_clk_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                     //  bfm_master_clk_reset_reset_bridge_in_reset.reset
		.jtag_master_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // jtag_master_clk_reset_reset_bridge_in_reset.reset
		.bfm_master_m0_address                             (bfm_master_m0_address),                              //                               bfm_master_m0.address
		.bfm_master_m0_waitrequest                         (bfm_master_m0_waitrequest),                          //                                            .waitrequest
		.bfm_master_m0_byteenable                          (bfm_master_m0_byteenable),                           //                                            .byteenable
		.bfm_master_m0_read                                (bfm_master_m0_read),                                 //                                            .read
		.bfm_master_m0_readdata                            (bfm_master_m0_readdata),                             //                                            .readdata
		.bfm_master_m0_readdatavalid                       (bfm_master_m0_readdatavalid),                        //                                            .readdatavalid
		.bfm_master_m0_write                               (bfm_master_m0_write),                                //                                            .write
		.bfm_master_m0_writedata                           (bfm_master_m0_writedata),                            //                                            .writedata
		.jtag_master_master_address                        (jtag_master_master_address),                         //                          jtag_master_master.address
		.jtag_master_master_waitrequest                    (jtag_master_master_waitrequest),                     //                                            .waitrequest
		.jtag_master_master_byteenable                     (jtag_master_master_byteenable),                      //                                            .byteenable
		.jtag_master_master_read                           (jtag_master_master_read),                            //                                            .read
		.jtag_master_master_readdata                       (jtag_master_master_readdata),                        //                                            .readdata
		.jtag_master_master_readdatavalid                  (jtag_master_master_readdatavalid),                   //                                            .readdatavalid
		.jtag_master_master_write                          (jtag_master_master_write),                           //                                            .write
		.jtag_master_master_writedata                      (jtag_master_master_writedata),                       //                                            .writedata
		.control_bits_s1_address                           (mm_interconnect_0_control_bits_s1_address),          //                             control_bits_s1.address
		.control_bits_s1_write                             (mm_interconnect_0_control_bits_s1_write),            //                                            .write
		.control_bits_s1_readdata                          (mm_interconnect_0_control_bits_s1_readdata),         //                                            .readdata
		.control_bits_s1_writedata                         (mm_interconnect_0_control_bits_s1_writedata),        //                                            .writedata
		.control_bits_s1_chipselect                        (mm_interconnect_0_control_bits_s1_chipselect),       //                                            .chipselect
		.dac_div_s1_address                                (mm_interconnect_0_dac_div_s1_address),               //                                  dac_div_s1.address
		.dac_div_s1_write                                  (mm_interconnect_0_dac_div_s1_write),                 //                                            .write
		.dac_div_s1_readdata                               (mm_interconnect_0_dac_div_s1_readdata),              //                                            .readdata
		.dac_div_s1_writedata                              (mm_interconnect_0_dac_div_s1_writedata),             //                                            .writedata
		.dac_div_s1_chipselect                             (mm_interconnect_0_dac_div_s1_chipselect),            //                                            .chipselect
		.dac_gain_s1_address                               (mm_interconnect_0_dac_gain_s1_address),              //                                 dac_gain_s1.address
		.dac_gain_s1_write                                 (mm_interconnect_0_dac_gain_s1_write),                //                                            .write
		.dac_gain_s1_readdata                              (mm_interconnect_0_dac_gain_s1_readdata),             //                                            .readdata
		.dac_gain_s1_writedata                             (mm_interconnect_0_dac_gain_s1_writedata),            //                                            .writedata
		.dac_gain_s1_chipselect                            (mm_interconnect_0_dac_gain_s1_chipselect),           //                                            .chipselect
		.gain_controller_s1_address                        (mm_interconnect_0_gain_controller_s1_address),       //                          gain_controller_s1.address
		.gain_controller_s1_write                          (mm_interconnect_0_gain_controller_s1_write),         //                                            .write
		.gain_controller_s1_readdata                       (mm_interconnect_0_gain_controller_s1_readdata),      //                                            .readdata
		.gain_controller_s1_writedata                      (mm_interconnect_0_gain_controller_s1_writedata),     //                                            .writedata
		.gain_controller_s1_chipselect                     (mm_interconnect_0_gain_controller_s1_chipselect),    //                                            .chipselect
		.lia_1_x_s1_address                                (mm_interconnect_0_lia_1_x_s1_address),               //                                  lia_1_x_s1.address
		.lia_1_x_s1_readdata                               (mm_interconnect_0_lia_1_x_s1_readdata),              //                                            .readdata
		.lia_1_y_s1_address                                (mm_interconnect_0_lia_1_y_s1_address),               //                                  lia_1_y_s1.address
		.lia_1_y_s1_readdata                               (mm_interconnect_0_lia_1_y_s1_readdata),              //                                            .readdata
		.nco_freq_control_1_s1_address                     (mm_interconnect_0_nco_freq_control_1_s1_address),    //                       nco_freq_control_1_s1.address
		.nco_freq_control_1_s1_write                       (mm_interconnect_0_nco_freq_control_1_s1_write),      //                                            .write
		.nco_freq_control_1_s1_readdata                    (mm_interconnect_0_nco_freq_control_1_s1_readdata),   //                                            .readdata
		.nco_freq_control_1_s1_writedata                   (mm_interconnect_0_nco_freq_control_1_s1_writedata),  //                                            .writedata
		.nco_freq_control_1_s1_chipselect                  (mm_interconnect_0_nco_freq_control_1_s1_chipselect), //                                            .chipselect
		.nco_freq_control_2_s1_address                     (mm_interconnect_0_nco_freq_control_2_s1_address),    //                       nco_freq_control_2_s1.address
		.nco_freq_control_2_s1_write                       (mm_interconnect_0_nco_freq_control_2_s1_write),      //                                            .write
		.nco_freq_control_2_s1_readdata                    (mm_interconnect_0_nco_freq_control_2_s1_readdata),   //                                            .readdata
		.nco_freq_control_2_s1_writedata                   (mm_interconnect_0_nco_freq_control_2_s1_writedata),  //                                            .writedata
		.nco_freq_control_2_s1_chipselect                  (mm_interconnect_0_nco_freq_control_2_s1_chipselect), //                                            .chipselect
		.nco_freq_ctrl_3_s1_address                        (mm_interconnect_0_nco_freq_ctrl_3_s1_address),       //                          nco_freq_ctrl_3_s1.address
		.nco_freq_ctrl_3_s1_write                          (mm_interconnect_0_nco_freq_ctrl_3_s1_write),         //                                            .write
		.nco_freq_ctrl_3_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_3_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_3_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_3_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_3_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect),    //                                            .chipselect
		.nco_freq_ctrl_4_s1_address                        (mm_interconnect_0_nco_freq_ctrl_4_s1_address),       //                          nco_freq_ctrl_4_s1.address
		.nco_freq_ctrl_4_s1_write                          (mm_interconnect_0_nco_freq_ctrl_4_s1_write),         //                                            .write
		.nco_freq_ctrl_4_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_4_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_4_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_4_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_4_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect),    //                                            .chipselect
		.nco_freq_ctrl_5_s1_address                        (mm_interconnect_0_nco_freq_ctrl_5_s1_address),       //                          nco_freq_ctrl_5_s1.address
		.nco_freq_ctrl_5_s1_write                          (mm_interconnect_0_nco_freq_ctrl_5_s1_write),         //                                            .write
		.nco_freq_ctrl_5_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_5_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_5_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_5_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_5_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect),    //                                            .chipselect
		.nco_freq_ctrl_6_s1_address                        (mm_interconnect_0_nco_freq_ctrl_6_s1_address),       //                          nco_freq_ctrl_6_s1.address
		.nco_freq_ctrl_6_s1_write                          (mm_interconnect_0_nco_freq_ctrl_6_s1_write),         //                                            .write
		.nco_freq_ctrl_6_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_6_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_6_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_6_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_6_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect),    //                                            .chipselect
		.nco_freq_ctrl_7_s1_address                        (mm_interconnect_0_nco_freq_ctrl_7_s1_address),       //                          nco_freq_ctrl_7_s1.address
		.nco_freq_ctrl_7_s1_write                          (mm_interconnect_0_nco_freq_ctrl_7_s1_write),         //                                            .write
		.nco_freq_ctrl_7_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_7_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_7_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_7_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_7_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect),    //                                            .chipselect
		.nco_freq_ctrl_8_s1_address                        (mm_interconnect_0_nco_freq_ctrl_8_s1_address),       //                          nco_freq_ctrl_8_s1.address
		.nco_freq_ctrl_8_s1_write                          (mm_interconnect_0_nco_freq_ctrl_8_s1_write),         //                                            .write
		.nco_freq_ctrl_8_s1_readdata                       (mm_interconnect_0_nco_freq_ctrl_8_s1_readdata),      //                                            .readdata
		.nco_freq_ctrl_8_s1_writedata                      (mm_interconnect_0_nco_freq_ctrl_8_s1_writedata),     //                                            .writedata
		.nco_freq_ctrl_8_s1_chipselect                     (mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect),    //                                            .chipselect
		.nco_phase_ctrl_1_s1_address                       (mm_interconnect_0_nco_phase_ctrl_1_s1_address),      //                         nco_phase_ctrl_1_s1.address
		.nco_phase_ctrl_1_s1_write                         (mm_interconnect_0_nco_phase_ctrl_1_s1_write),        //                                            .write
		.nco_phase_ctrl_1_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_1_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_1_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_1_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_1_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_2_s1_address                       (mm_interconnect_0_nco_phase_ctrl_2_s1_address),      //                         nco_phase_ctrl_2_s1.address
		.nco_phase_ctrl_2_s1_write                         (mm_interconnect_0_nco_phase_ctrl_2_s1_write),        //                                            .write
		.nco_phase_ctrl_2_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_2_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_2_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_2_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_2_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_3_s1_address                       (mm_interconnect_0_nco_phase_ctrl_3_s1_address),      //                         nco_phase_ctrl_3_s1.address
		.nco_phase_ctrl_3_s1_write                         (mm_interconnect_0_nco_phase_ctrl_3_s1_write),        //                                            .write
		.nco_phase_ctrl_3_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_3_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_3_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_3_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_3_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_4_s1_address                       (mm_interconnect_0_nco_phase_ctrl_4_s1_address),      //                         nco_phase_ctrl_4_s1.address
		.nco_phase_ctrl_4_s1_write                         (mm_interconnect_0_nco_phase_ctrl_4_s1_write),        //                                            .write
		.nco_phase_ctrl_4_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_4_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_4_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_4_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_4_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_5_s1_address                       (mm_interconnect_0_nco_phase_ctrl_5_s1_address),      //                         nco_phase_ctrl_5_s1.address
		.nco_phase_ctrl_5_s1_write                         (mm_interconnect_0_nco_phase_ctrl_5_s1_write),        //                                            .write
		.nco_phase_ctrl_5_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_5_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_5_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_5_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_5_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_6_s1_address                       (mm_interconnect_0_nco_phase_ctrl_6_s1_address),      //                         nco_phase_ctrl_6_s1.address
		.nco_phase_ctrl_6_s1_write                         (mm_interconnect_0_nco_phase_ctrl_6_s1_write),        //                                            .write
		.nco_phase_ctrl_6_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_6_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_6_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_6_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_6_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_7_s1_address                       (mm_interconnect_0_nco_phase_ctrl_7_s1_address),      //                         nco_phase_ctrl_7_s1.address
		.nco_phase_ctrl_7_s1_write                         (mm_interconnect_0_nco_phase_ctrl_7_s1_write),        //                                            .write
		.nco_phase_ctrl_7_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_7_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_7_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_7_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_7_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect),   //                                            .chipselect
		.nco_phase_ctrl_8_s1_address                       (mm_interconnect_0_nco_phase_ctrl_8_s1_address),      //                         nco_phase_ctrl_8_s1.address
		.nco_phase_ctrl_8_s1_write                         (mm_interconnect_0_nco_phase_ctrl_8_s1_write),        //                                            .write
		.nco_phase_ctrl_8_s1_readdata                      (mm_interconnect_0_nco_phase_ctrl_8_s1_readdata),     //                                            .readdata
		.nco_phase_ctrl_8_s1_writedata                     (mm_interconnect_0_nco_phase_ctrl_8_s1_writedata),    //                                            .writedata
		.nco_phase_ctrl_8_s1_chipselect                    (mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect),   //                                            .chipselect
		.onchip_ram_s1_address                             (mm_interconnect_0_onchip_ram_s1_address),            //                               onchip_ram_s1.address
		.onchip_ram_s1_write                               (mm_interconnect_0_onchip_ram_s1_write),              //                                            .write
		.onchip_ram_s1_readdata                            (mm_interconnect_0_onchip_ram_s1_readdata),           //                                            .readdata
		.onchip_ram_s1_writedata                           (mm_interconnect_0_onchip_ram_s1_writedata),          //                                            .writedata
		.onchip_ram_s1_byteenable                          (mm_interconnect_0_onchip_ram_s1_byteenable),         //                                            .byteenable
		.onchip_ram_s1_chipselect                          (mm_interconnect_0_onchip_ram_s1_chipselect),         //                                            .chipselect
		.onchip_ram_s1_clken                               (mm_interconnect_0_onchip_ram_s1_clken)               //                                            .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
