-- qsys_system.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qsys_system is
	port (
		clk_clk             : in  std_logic                     := '0'; --          clk.clk
		gain_ctrl_export    : out std_logic_vector(5 downto 0);         --    gain_ctrl.export
		phase_incr_1_export : out std_logic_vector(19 downto 0);        -- phase_incr_1.export
		phase_incr_2_export : out std_logic_vector(19 downto 0);        -- phase_incr_2.export
		phase_incr_3_export : out std_logic_vector(19 downto 0);        -- phase_incr_3.export
		phase_incr_4_export : out std_logic_vector(19 downto 0);        -- phase_incr_4.export
		phase_incr_5_export : out std_logic_vector(19 downto 0);        -- phase_incr_5.export
		phase_incr_6_export : out std_logic_vector(19 downto 0);        -- phase_incr_6.export
		phase_incr_7_export : out std_logic_vector(19 downto 0);        -- phase_incr_7.export
		phase_incr_8_export : out std_logic_vector(19 downto 0);        -- phase_incr_8.export
		phase_offs_1_export : out std_logic_vector(19 downto 0);        -- phase_offs_1.export
		phase_offs_2_export : out std_logic_vector(19 downto 0);        -- phase_offs_2.export
		phase_offs_3_export : out std_logic_vector(19 downto 0);        -- phase_offs_3.export
		phase_offs_4_export : out std_logic_vector(19 downto 0);        -- phase_offs_4.export
		phase_offs_5_export : out std_logic_vector(19 downto 0);        -- phase_offs_5.export
		phase_offs_6_export : out std_logic_vector(19 downto 0);        -- phase_offs_6.export
		phase_offs_7_export : out std_logic_vector(19 downto 0);        -- phase_offs_7.export
		phase_offs_8_export : out std_logic_vector(19 downto 0);        -- phase_offs_8.export
		reset_reset_n       : in  std_logic                     := '0'; --        reset.reset_n
		resetrequest_reset  : out std_logic                             -- resetrequest.reset
	);
end entity qsys_system;

architecture rtl of qsys_system is
	component altera_avalon_mm_master_bfm is
		generic (
			AV_ADDRESS_W               : integer := 32;
			AV_SYMBOL_W                : integer := 8;
			AV_NUMSYMBOLS              : integer := 4;
			AV_BURSTCOUNT_W            : integer := 3;
			AV_READRESPONSE_W          : integer := 8;
			AV_WRITERESPONSE_W         : integer := 8;
			USE_READ                   : integer := 1;
			USE_WRITE                  : integer := 1;
			USE_ADDRESS                : integer := 1;
			USE_BYTE_ENABLE            : integer := 1;
			USE_BURSTCOUNT             : integer := 1;
			USE_READ_DATA              : integer := 1;
			USE_READ_DATA_VALID        : integer := 1;
			USE_WRITE_DATA             : integer := 1;
			USE_BEGIN_TRANSFER         : integer := 0;
			USE_BEGIN_BURST_TRANSFER   : integer := 0;
			USE_WAIT_REQUEST           : integer := 1;
			USE_TRANSACTIONID          : integer := 0;
			USE_WRITERESPONSE          : integer := 0;
			USE_READRESPONSE           : integer := 0;
			USE_CLKEN                  : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR : integer := 1;
			AV_BURST_LINEWRAP          : integer := 1;
			AV_BURST_BNDR_ONLY         : integer := 1;
			AV_MAX_PENDING_READS       : integer := 0;
			AV_MAX_PENDING_WRITES      : integer := 0;
			AV_FIX_READ_LATENCY        : integer := 1;
			AV_READ_WAIT_TIME          : integer := 1;
			AV_WRITE_WAIT_TIME         : integer := 0;
			REGISTER_WAITREQUEST       : integer := 0;
			AV_REGISTERINCOMINGSIGNALS : integer := 0;
			VHDL_ID                    : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			avm_address            : out std_logic_vector(31 downto 0);                    -- address
			avm_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			avm_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			avm_write              : out std_logic;                                        -- write
			avm_read               : out std_logic;                                        -- read
			avm_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			avm_burstcount         : out std_logic_vector(2 downto 0);                     -- burstcount
			avm_begintransfer      : out std_logic;                                        -- begintransfer
			avm_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			avm_arbiterlock        : out std_logic;                                        -- arbiterlock
			avm_lock               : out std_logic;                                        -- lock
			avm_debugaccess        : out std_logic;                                        -- debugaccess
			avm_transactionid      : out std_logic_vector(7 downto 0);                     -- transactionid
			avm_readid             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readid
			avm_writeid            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writeid
			avm_clken              : out std_logic;                                        -- clken
			avm_response           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			avm_writeresponsevalid : in  std_logic                     := 'X';             -- writeresponsevalid
			avm_readresponse       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readresponse
			avm_writeresponse      : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- writeresponse
		);
	end component altera_avalon_mm_master_bfm;

	component qsys_system_gain_controller is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component qsys_system_gain_controller;

	component qsys_system_jtag_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component qsys_system_jtag_master;

	component qsys_system_nco_freq_control_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(19 downto 0)                     -- export
		);
	end component qsys_system_nco_freq_control_1;

	component qsys_system_nco_freq_control_2 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(19 downto 0)                     -- export
		);
	end component qsys_system_nco_freq_control_2;

	component qsys_system_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component qsys_system_onchip_ram;

	component qsys_system_mm_interconnect_0 is
		port (
			clk_clk_clk                                       : in  std_logic                     := 'X';             -- clk
			bfm_master_clk_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			jtag_master_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			bfm_master_m0_address                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			bfm_master_m0_waitrequest                         : out std_logic;                                        -- waitrequest
			bfm_master_m0_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			bfm_master_m0_read                                : in  std_logic                     := 'X';             -- read
			bfm_master_m0_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			bfm_master_m0_readdatavalid                       : out std_logic;                                        -- readdatavalid
			bfm_master_m0_write                               : in  std_logic                     := 'X';             -- write
			bfm_master_m0_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			jtag_master_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			jtag_master_master_waitrequest                    : out std_logic;                                        -- waitrequest
			jtag_master_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_master_master_read                           : in  std_logic                     := 'X';             -- read
			jtag_master_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_master_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			jtag_master_master_write                          : in  std_logic                     := 'X';             -- write
			jtag_master_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			gain_controller_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			gain_controller_s1_write                          : out std_logic;                                        -- write
			gain_controller_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			gain_controller_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			gain_controller_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_control_1_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_control_1_s1_write                       : out std_logic;                                        -- write
			nco_freq_control_1_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_control_1_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_control_1_s1_chipselect                  : out std_logic;                                        -- chipselect
			nco_freq_control_2_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_control_2_s1_write                       : out std_logic;                                        -- write
			nco_freq_control_2_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_control_2_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_control_2_s1_chipselect                  : out std_logic;                                        -- chipselect
			nco_freq_ctrl_3_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_3_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_3_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_3_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_3_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_ctrl_4_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_4_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_4_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_4_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_4_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_ctrl_5_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_5_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_5_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_5_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_5_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_ctrl_6_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_6_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_6_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_6_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_6_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_ctrl_7_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_7_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_7_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_7_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_7_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_freq_ctrl_8_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			nco_freq_ctrl_8_s1_write                          : out std_logic;                                        -- write
			nco_freq_ctrl_8_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_freq_ctrl_8_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			nco_freq_ctrl_8_s1_chipselect                     : out std_logic;                                        -- chipselect
			nco_phase_ctrl_1_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_1_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_1_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_1_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_1_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_2_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_2_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_2_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_2_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_2_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_3_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_3_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_3_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_3_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_3_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_4_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_4_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_4_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_4_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_4_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_5_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_5_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_5_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_5_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_5_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_6_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_6_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_6_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_6_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_6_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_7_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_7_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_7_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_7_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_7_s1_chipselect                    : out std_logic;                                        -- chipselect
			nco_phase_ctrl_8_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			nco_phase_ctrl_8_s1_write                         : out std_logic;                                        -- write
			nco_phase_ctrl_8_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nco_phase_ctrl_8_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			nco_phase_ctrl_8_s1_chipselect                    : out std_logic;                                        -- chipselect
			onchip_ram_s1_address                             : out std_logic_vector(9 downto 0);                     -- address
			onchip_ram_s1_write                               : out std_logic;                                        -- write
			onchip_ram_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                          : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                               : out std_logic                                         -- clken
		);
	end component qsys_system_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal bfm_master_m0_readdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:bfm_master_m0_readdata -> bfm_master:avm_readdata
	signal bfm_master_m0_waitrequest                               : std_logic;                     -- mm_interconnect_0:bfm_master_m0_waitrequest -> bfm_master:avm_waitrequest
	signal bfm_master_m0_address                                   : std_logic_vector(31 downto 0); -- bfm_master:avm_address -> mm_interconnect_0:bfm_master_m0_address
	signal bfm_master_m0_read                                      : std_logic;                     -- bfm_master:avm_read -> mm_interconnect_0:bfm_master_m0_read
	signal bfm_master_m0_byteenable                                : std_logic_vector(3 downto 0);  -- bfm_master:avm_byteenable -> mm_interconnect_0:bfm_master_m0_byteenable
	signal bfm_master_m0_readdatavalid                             : std_logic;                     -- mm_interconnect_0:bfm_master_m0_readdatavalid -> bfm_master:avm_readdatavalid
	signal bfm_master_m0_writedata                                 : std_logic_vector(31 downto 0); -- bfm_master:avm_writedata -> mm_interconnect_0:bfm_master_m0_writedata
	signal bfm_master_m0_write                                     : std_logic;                     -- bfm_master:avm_write -> mm_interconnect_0:bfm_master_m0_write
	signal jtag_master_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	signal jtag_master_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	signal jtag_master_master_address                              : std_logic_vector(31 downto 0); -- jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	signal jtag_master_master_read                                 : std_logic;                     -- jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	signal jtag_master_master_byteenable                           : std_logic_vector(3 downto 0);  -- jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	signal jtag_master_master_readdatavalid                        : std_logic;                     -- mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	signal jtag_master_master_write                                : std_logic;                     -- jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	signal jtag_master_master_writedata                            : std_logic_vector(31 downto 0); -- jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	signal mm_interconnect_0_nco_freq_control_1_s1_chipselect      : std_logic;                     -- mm_interconnect_0:nco_freq_control_1_s1_chipselect -> nco_freq_control_1:chipselect
	signal mm_interconnect_0_nco_freq_control_1_s1_readdata        : std_logic_vector(31 downto 0); -- nco_freq_control_1:readdata -> mm_interconnect_0:nco_freq_control_1_s1_readdata
	signal mm_interconnect_0_nco_freq_control_1_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_control_1_s1_address -> nco_freq_control_1:address
	signal mm_interconnect_0_nco_freq_control_1_s1_write           : std_logic;                     -- mm_interconnect_0:nco_freq_control_1_s1_write -> mm_interconnect_0_nco_freq_control_1_s1_write:in
	signal mm_interconnect_0_nco_freq_control_1_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_control_1_s1_writedata -> nco_freq_control_1:writedata
	signal mm_interconnect_0_nco_freq_control_2_s1_chipselect      : std_logic;                     -- mm_interconnect_0:nco_freq_control_2_s1_chipselect -> nco_freq_control_2:chipselect
	signal mm_interconnect_0_nco_freq_control_2_s1_readdata        : std_logic_vector(31 downto 0); -- nco_freq_control_2:readdata -> mm_interconnect_0:nco_freq_control_2_s1_readdata
	signal mm_interconnect_0_nco_freq_control_2_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_control_2_s1_address -> nco_freq_control_2:address
	signal mm_interconnect_0_nco_freq_control_2_s1_write           : std_logic;                     -- mm_interconnect_0:nco_freq_control_2_s1_write -> mm_interconnect_0_nco_freq_control_2_s1_write:in
	signal mm_interconnect_0_nco_freq_control_2_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_control_2_s1_writedata -> nco_freq_control_2:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect              : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                 : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                   : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                   : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_1_s1_chipselect -> nco_phase_ctrl_1:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_1:readdata -> mm_interconnect_0:nco_phase_ctrl_1_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_1_s1_address -> nco_phase_ctrl_1:address
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_1_s1_write -> mm_interconnect_0_nco_phase_ctrl_1_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_1_s1_writedata -> nco_phase_ctrl_1:writedata
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_2_s1_chipselect -> nco_phase_ctrl_2:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_2:readdata -> mm_interconnect_0:nco_phase_ctrl_2_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_2_s1_address -> nco_phase_ctrl_2:address
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_2_s1_write -> mm_interconnect_0_nco_phase_ctrl_2_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_2_s1_writedata -> nco_phase_ctrl_2:writedata
	signal mm_interconnect_0_gain_controller_s1_chipselect         : std_logic;                     -- mm_interconnect_0:gain_controller_s1_chipselect -> gain_controller:chipselect
	signal mm_interconnect_0_gain_controller_s1_readdata           : std_logic_vector(31 downto 0); -- gain_controller:readdata -> mm_interconnect_0:gain_controller_s1_readdata
	signal mm_interconnect_0_gain_controller_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:gain_controller_s1_address -> gain_controller:address
	signal mm_interconnect_0_gain_controller_s1_write              : std_logic;                     -- mm_interconnect_0:gain_controller_s1_write -> mm_interconnect_0_gain_controller_s1_write:in
	signal mm_interconnect_0_gain_controller_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:gain_controller_s1_writedata -> gain_controller:writedata
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_3_s1_chipselect -> nco_freq_ctrl_3:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_3:readdata -> mm_interconnect_0:nco_freq_ctrl_3_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_3_s1_address -> nco_freq_ctrl_3:address
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_3_s1_write -> mm_interconnect_0_nco_freq_ctrl_3_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_3_s1_writedata -> nco_freq_ctrl_3:writedata
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_4_s1_chipselect -> nco_freq_ctrl_4:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_4:readdata -> mm_interconnect_0:nco_freq_ctrl_4_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_4_s1_address -> nco_freq_ctrl_4:address
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_4_s1_write -> mm_interconnect_0_nco_freq_ctrl_4_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_4_s1_writedata -> nco_freq_ctrl_4:writedata
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_5_s1_chipselect -> nco_freq_ctrl_5:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_5:readdata -> mm_interconnect_0:nco_freq_ctrl_5_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_5_s1_address -> nco_freq_ctrl_5:address
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_5_s1_write -> mm_interconnect_0_nco_freq_ctrl_5_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_5_s1_writedata -> nco_freq_ctrl_5:writedata
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_6_s1_chipselect -> nco_freq_ctrl_6:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_6:readdata -> mm_interconnect_0:nco_freq_ctrl_6_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_6_s1_address -> nco_freq_ctrl_6:address
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_6_s1_write -> mm_interconnect_0_nco_freq_ctrl_6_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_6_s1_writedata -> nco_freq_ctrl_6:writedata
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_7_s1_chipselect -> nco_freq_ctrl_7:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_7:readdata -> mm_interconnect_0:nco_freq_ctrl_7_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_7_s1_address -> nco_freq_ctrl_7:address
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_7_s1_write -> mm_interconnect_0_nco_freq_ctrl_7_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_7_s1_writedata -> nco_freq_ctrl_7:writedata
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect         : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_8_s1_chipselect -> nco_freq_ctrl_8:chipselect
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_readdata           : std_logic_vector(31 downto 0); -- nco_freq_ctrl_8:readdata -> mm_interconnect_0:nco_freq_ctrl_8_s1_readdata
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_freq_ctrl_8_s1_address -> nco_freq_ctrl_8:address
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_write              : std_logic;                     -- mm_interconnect_0:nco_freq_ctrl_8_s1_write -> mm_interconnect_0_nco_freq_ctrl_8_s1_write:in
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_freq_ctrl_8_s1_writedata -> nco_freq_ctrl_8:writedata
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_3_s1_chipselect -> nco_phase_ctrl_3:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_3:readdata -> mm_interconnect_0:nco_phase_ctrl_3_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_3_s1_address -> nco_phase_ctrl_3:address
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_3_s1_write -> mm_interconnect_0_nco_phase_ctrl_3_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_3_s1_writedata -> nco_phase_ctrl_3:writedata
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_4_s1_chipselect -> nco_phase_ctrl_4:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_4:readdata -> mm_interconnect_0:nco_phase_ctrl_4_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_4_s1_address -> nco_phase_ctrl_4:address
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_4_s1_write -> mm_interconnect_0_nco_phase_ctrl_4_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_4_s1_writedata -> nco_phase_ctrl_4:writedata
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_5_s1_chipselect -> nco_phase_ctrl_5:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_5:readdata -> mm_interconnect_0:nco_phase_ctrl_5_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_5_s1_address -> nco_phase_ctrl_5:address
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_5_s1_write -> mm_interconnect_0_nco_phase_ctrl_5_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_5_s1_writedata -> nco_phase_ctrl_5:writedata
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_6_s1_chipselect -> nco_phase_ctrl_6:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_6:readdata -> mm_interconnect_0:nco_phase_ctrl_6_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_6_s1_address -> nco_phase_ctrl_6:address
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_6_s1_write -> mm_interconnect_0_nco_phase_ctrl_6_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_6_s1_writedata -> nco_phase_ctrl_6:writedata
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_7_s1_chipselect -> nco_phase_ctrl_7:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_7:readdata -> mm_interconnect_0:nco_phase_ctrl_7_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_7_s1_address -> nco_phase_ctrl_7:address
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_7_s1_write -> mm_interconnect_0_nco_phase_ctrl_7_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_7_s1_writedata -> nco_phase_ctrl_7:writedata
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect        : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_8_s1_chipselect -> nco_phase_ctrl_8:chipselect
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_readdata          : std_logic_vector(31 downto 0); -- nco_phase_ctrl_8:readdata -> mm_interconnect_0:nco_phase_ctrl_8_s1_readdata
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_address           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:nco_phase_ctrl_8_s1_address -> nco_phase_ctrl_8:address
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_write             : std_logic;                     -- mm_interconnect_0:nco_phase_ctrl_8_s1_write -> mm_interconnect_0_nco_phase_ctrl_8_s1_write:in
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:nco_phase_ctrl_8_s1_writedata -> nco_phase_ctrl_8:writedata
	signal rst_controller_reset_out_reset                          : std_logic;                     -- rst_controller:reset_out -> [bfm_master:reset, mm_interconnect_0:bfm_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                      : std_logic;                     -- rst_controller:reset_req -> [onchip_ram:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                 : std_logic;                     -- reset_reset_n:inv -> [jtag_master:clk_reset_reset, rst_controller:reset_in0]
	signal mm_interconnect_0_nco_freq_control_1_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_nco_freq_control_1_s1_write:inv -> nco_freq_control_1:write_n
	signal mm_interconnect_0_nco_freq_control_2_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_nco_freq_control_2_s1_write:inv -> nco_freq_control_2:write_n
	signal mm_interconnect_0_nco_phase_ctrl_1_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_1_s1_write:inv -> nco_phase_ctrl_1:write_n
	signal mm_interconnect_0_nco_phase_ctrl_2_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_2_s1_write:inv -> nco_phase_ctrl_2:write_n
	signal mm_interconnect_0_gain_controller_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_gain_controller_s1_write:inv -> gain_controller:write_n
	signal mm_interconnect_0_nco_freq_ctrl_3_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_3_s1_write:inv -> nco_freq_ctrl_3:write_n
	signal mm_interconnect_0_nco_freq_ctrl_4_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_4_s1_write:inv -> nco_freq_ctrl_4:write_n
	signal mm_interconnect_0_nco_freq_ctrl_5_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_5_s1_write:inv -> nco_freq_ctrl_5:write_n
	signal mm_interconnect_0_nco_freq_ctrl_6_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_6_s1_write:inv -> nco_freq_ctrl_6:write_n
	signal mm_interconnect_0_nco_freq_ctrl_7_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_7_s1_write:inv -> nco_freq_ctrl_7:write_n
	signal mm_interconnect_0_nco_freq_ctrl_8_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_nco_freq_ctrl_8_s1_write:inv -> nco_freq_ctrl_8:write_n
	signal mm_interconnect_0_nco_phase_ctrl_3_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_3_s1_write:inv -> nco_phase_ctrl_3:write_n
	signal mm_interconnect_0_nco_phase_ctrl_4_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_4_s1_write:inv -> nco_phase_ctrl_4:write_n
	signal mm_interconnect_0_nco_phase_ctrl_5_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_5_s1_write:inv -> nco_phase_ctrl_5:write_n
	signal mm_interconnect_0_nco_phase_ctrl_6_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_6_s1_write:inv -> nco_phase_ctrl_6:write_n
	signal mm_interconnect_0_nco_phase_ctrl_7_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_7_s1_write:inv -> nco_phase_ctrl_7:write_n
	signal mm_interconnect_0_nco_phase_ctrl_8_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_nco_phase_ctrl_8_s1_write:inv -> nco_phase_ctrl_8:write_n
	signal rst_controller_reset_out_reset_ports_inv                : std_logic;                     -- rst_controller_reset_out_reset:inv -> [gain_controller:reset_n, nco_freq_control_1:reset_n, nco_freq_control_2:reset_n, nco_freq_ctrl_3:reset_n, nco_freq_ctrl_4:reset_n, nco_freq_ctrl_5:reset_n, nco_freq_ctrl_6:reset_n, nco_freq_ctrl_7:reset_n, nco_freq_ctrl_8:reset_n, nco_phase_ctrl_1:reset_n, nco_phase_ctrl_2:reset_n, nco_phase_ctrl_3:reset_n, nco_phase_ctrl_4:reset_n, nco_phase_ctrl_5:reset_n, nco_phase_ctrl_6:reset_n, nco_phase_ctrl_7:reset_n, nco_phase_ctrl_8:reset_n]

begin

	bfm_master : component altera_avalon_mm_master_bfm
		generic map (
			AV_ADDRESS_W               => 32,
			AV_SYMBOL_W                => 8,
			AV_NUMSYMBOLS              => 4,
			AV_BURSTCOUNT_W            => 3,
			AV_READRESPONSE_W          => 8,
			AV_WRITERESPONSE_W         => 8,
			USE_READ                   => 1,
			USE_WRITE                  => 1,
			USE_ADDRESS                => 1,
			USE_BYTE_ENABLE            => 1,
			USE_BURSTCOUNT             => 0,
			USE_READ_DATA              => 1,
			USE_READ_DATA_VALID        => 1,
			USE_WRITE_DATA             => 1,
			USE_BEGIN_TRANSFER         => 0,
			USE_BEGIN_BURST_TRANSFER   => 0,
			USE_WAIT_REQUEST           => 1,
			USE_TRANSACTIONID          => 0,
			USE_WRITERESPONSE          => 0,
			USE_READRESPONSE           => 0,
			USE_CLKEN                  => 0,
			AV_CONSTANT_BURST_BEHAVIOR => 1,
			AV_BURST_LINEWRAP          => 1,
			AV_BURST_BNDR_ONLY         => 1,
			AV_MAX_PENDING_READS       => 0,
			AV_MAX_PENDING_WRITES      => 0,
			AV_FIX_READ_LATENCY        => 1,
			AV_READ_WAIT_TIME          => 1,
			AV_WRITE_WAIT_TIME         => 0,
			REGISTER_WAITREQUEST       => 0,
			AV_REGISTERINCOMINGSIGNALS => 0,
			VHDL_ID                    => 0
		)
		port map (
			clk                    => clk_clk,                        --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			avm_address            => bfm_master_m0_address,          --        m0.address
			avm_readdata           => bfm_master_m0_readdata,         --          .readdata
			avm_writedata          => bfm_master_m0_writedata,        --          .writedata
			avm_waitrequest        => bfm_master_m0_waitrequest,      --          .waitrequest
			avm_write              => bfm_master_m0_write,            --          .write
			avm_read               => bfm_master_m0_read,             --          .read
			avm_byteenable         => bfm_master_m0_byteenable,       --          .byteenable
			avm_readdatavalid      => bfm_master_m0_readdatavalid,    --          .readdatavalid
			avm_burstcount         => open,                           -- (terminated)
			avm_begintransfer      => open,                           -- (terminated)
			avm_beginbursttransfer => open,                           -- (terminated)
			avm_arbiterlock        => open,                           -- (terminated)
			avm_lock               => open,                           -- (terminated)
			avm_debugaccess        => open,                           -- (terminated)
			avm_transactionid      => open,                           -- (terminated)
			avm_readid             => "00000000",                     -- (terminated)
			avm_writeid            => "00000000",                     -- (terminated)
			avm_clken              => open,                           -- (terminated)
			avm_response           => "00",                           -- (terminated)
			avm_writeresponsevalid => '0',                            -- (terminated)
			avm_readresponse       => "00000000",                     -- (terminated)
			avm_writeresponse      => "00000000"                      -- (terminated)
		);

	gain_controller : component qsys_system_gain_controller
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_gain_controller_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_gain_controller_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_gain_controller_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_gain_controller_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_gain_controller_s1_readdata,        --                    .readdata
			out_port   => gain_ctrl_export                                      -- external_connection.export
		);

	jtag_master : component qsys_system_jtag_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                          --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,          --    clk_reset.reset
			master_address       => jtag_master_master_address,       --       master.address
			master_readdata      => jtag_master_master_readdata,      --             .readdata
			master_read          => jtag_master_master_read,          --             .read
			master_write         => jtag_master_master_write,         --             .write
			master_writedata     => jtag_master_master_writedata,     --             .writedata
			master_waitrequest   => jtag_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_master_master_byteenable,    --             .byteenable
			master_reset_reset   => resetrequest_reset                -- master_reset.reset
		);

	nco_freq_control_1 : component qsys_system_nco_freq_control_1
		port map (
			clk        => clk_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_control_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_control_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_control_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_control_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_control_1_s1_readdata,        --                    .readdata
			out_port   => phase_incr_1_export                                      -- external_connection.export
		);

	nco_freq_control_2 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_control_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_control_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_control_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_control_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_control_2_s1_readdata,        --                    .readdata
			out_port   => phase_incr_2_export                                      -- external_connection.export
		);

	nco_freq_ctrl_3 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_3_s1_readdata,        --                    .readdata
			out_port   => phase_incr_3_export                                   -- external_connection.export
		);

	nco_freq_ctrl_4 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_4_s1_readdata,        --                    .readdata
			out_port   => phase_incr_4_export                                   -- external_connection.export
		);

	nco_freq_ctrl_5 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_5_s1_readdata,        --                    .readdata
			out_port   => phase_incr_5_export                                   -- external_connection.export
		);

	nco_freq_ctrl_6 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_6_s1_readdata,        --                    .readdata
			out_port   => phase_incr_6_export                                   -- external_connection.export
		);

	nco_freq_ctrl_7 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_7_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_7_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_7_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_7_s1_readdata,        --                    .readdata
			out_port   => phase_incr_7_export                                   -- external_connection.export
		);

	nco_freq_ctrl_8 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => mm_interconnect_0_nco_freq_ctrl_8_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_freq_ctrl_8_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_freq_ctrl_8_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_freq_ctrl_8_s1_readdata,        --                    .readdata
			out_port   => phase_incr_8_export                                   -- external_connection.export
		);

	nco_phase_ctrl_1 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_1_s1_readdata,        --                    .readdata
			out_port   => phase_offs_1_export                                    -- external_connection.export
		);

	nco_phase_ctrl_2 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_2_s1_readdata,        --                    .readdata
			out_port   => phase_offs_2_export                                    -- external_connection.export
		);

	nco_phase_ctrl_3 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_3_s1_readdata,        --                    .readdata
			out_port   => phase_offs_3_export                                    -- external_connection.export
		);

	nco_phase_ctrl_4 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_4_s1_readdata,        --                    .readdata
			out_port   => phase_offs_4_export                                    -- external_connection.export
		);

	nco_phase_ctrl_5 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_5_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_5_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_5_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_5_s1_readdata,        --                    .readdata
			out_port   => phase_offs_5_export                                    -- external_connection.export
		);

	nco_phase_ctrl_6 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_6_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_6_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_6_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_6_s1_readdata,        --                    .readdata
			out_port   => phase_offs_6_export                                    -- external_connection.export
		);

	nco_phase_ctrl_7 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_7_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_7_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_7_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_7_s1_readdata,        --                    .readdata
			out_port   => phase_offs_7_export                                    -- external_connection.export
		);

	nco_phase_ctrl_8 : component qsys_system_nco_freq_control_2
		port map (
			clk        => clk_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_nco_phase_ctrl_8_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_nco_phase_ctrl_8_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_nco_phase_ctrl_8_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_nco_phase_ctrl_8_s1_readdata,        --                    .readdata
			out_port   => phase_offs_8_export                                    -- external_connection.export
		);

	onchip_ram : component qsys_system_onchip_ram
		port map (
			clk        => clk_clk,                                    --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	mm_interconnect_0 : component qsys_system_mm_interconnect_0
		port map (
			clk_clk_clk                                       => clk_clk,                                            --                                     clk_clk.clk
			bfm_master_clk_reset_reset_bridge_in_reset_reset  => rst_controller_reset_out_reset,                     --  bfm_master_clk_reset_reset_bridge_in_reset.reset
			jtag_master_clk_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                     -- jtag_master_clk_reset_reset_bridge_in_reset.reset
			bfm_master_m0_address                             => bfm_master_m0_address,                              --                               bfm_master_m0.address
			bfm_master_m0_waitrequest                         => bfm_master_m0_waitrequest,                          --                                            .waitrequest
			bfm_master_m0_byteenable                          => bfm_master_m0_byteenable,                           --                                            .byteenable
			bfm_master_m0_read                                => bfm_master_m0_read,                                 --                                            .read
			bfm_master_m0_readdata                            => bfm_master_m0_readdata,                             --                                            .readdata
			bfm_master_m0_readdatavalid                       => bfm_master_m0_readdatavalid,                        --                                            .readdatavalid
			bfm_master_m0_write                               => bfm_master_m0_write,                                --                                            .write
			bfm_master_m0_writedata                           => bfm_master_m0_writedata,                            --                                            .writedata
			jtag_master_master_address                        => jtag_master_master_address,                         --                          jtag_master_master.address
			jtag_master_master_waitrequest                    => jtag_master_master_waitrequest,                     --                                            .waitrequest
			jtag_master_master_byteenable                     => jtag_master_master_byteenable,                      --                                            .byteenable
			jtag_master_master_read                           => jtag_master_master_read,                            --                                            .read
			jtag_master_master_readdata                       => jtag_master_master_readdata,                        --                                            .readdata
			jtag_master_master_readdatavalid                  => jtag_master_master_readdatavalid,                   --                                            .readdatavalid
			jtag_master_master_write                          => jtag_master_master_write,                           --                                            .write
			jtag_master_master_writedata                      => jtag_master_master_writedata,                       --                                            .writedata
			gain_controller_s1_address                        => mm_interconnect_0_gain_controller_s1_address,       --                          gain_controller_s1.address
			gain_controller_s1_write                          => mm_interconnect_0_gain_controller_s1_write,         --                                            .write
			gain_controller_s1_readdata                       => mm_interconnect_0_gain_controller_s1_readdata,      --                                            .readdata
			gain_controller_s1_writedata                      => mm_interconnect_0_gain_controller_s1_writedata,     --                                            .writedata
			gain_controller_s1_chipselect                     => mm_interconnect_0_gain_controller_s1_chipselect,    --                                            .chipselect
			nco_freq_control_1_s1_address                     => mm_interconnect_0_nco_freq_control_1_s1_address,    --                       nco_freq_control_1_s1.address
			nco_freq_control_1_s1_write                       => mm_interconnect_0_nco_freq_control_1_s1_write,      --                                            .write
			nco_freq_control_1_s1_readdata                    => mm_interconnect_0_nco_freq_control_1_s1_readdata,   --                                            .readdata
			nco_freq_control_1_s1_writedata                   => mm_interconnect_0_nco_freq_control_1_s1_writedata,  --                                            .writedata
			nco_freq_control_1_s1_chipselect                  => mm_interconnect_0_nco_freq_control_1_s1_chipselect, --                                            .chipselect
			nco_freq_control_2_s1_address                     => mm_interconnect_0_nco_freq_control_2_s1_address,    --                       nco_freq_control_2_s1.address
			nco_freq_control_2_s1_write                       => mm_interconnect_0_nco_freq_control_2_s1_write,      --                                            .write
			nco_freq_control_2_s1_readdata                    => mm_interconnect_0_nco_freq_control_2_s1_readdata,   --                                            .readdata
			nco_freq_control_2_s1_writedata                   => mm_interconnect_0_nco_freq_control_2_s1_writedata,  --                                            .writedata
			nco_freq_control_2_s1_chipselect                  => mm_interconnect_0_nco_freq_control_2_s1_chipselect, --                                            .chipselect
			nco_freq_ctrl_3_s1_address                        => mm_interconnect_0_nco_freq_ctrl_3_s1_address,       --                          nco_freq_ctrl_3_s1.address
			nco_freq_ctrl_3_s1_write                          => mm_interconnect_0_nco_freq_ctrl_3_s1_write,         --                                            .write
			nco_freq_ctrl_3_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_3_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_3_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_3_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_3_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_3_s1_chipselect,    --                                            .chipselect
			nco_freq_ctrl_4_s1_address                        => mm_interconnect_0_nco_freq_ctrl_4_s1_address,       --                          nco_freq_ctrl_4_s1.address
			nco_freq_ctrl_4_s1_write                          => mm_interconnect_0_nco_freq_ctrl_4_s1_write,         --                                            .write
			nco_freq_ctrl_4_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_4_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_4_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_4_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_4_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_4_s1_chipselect,    --                                            .chipselect
			nco_freq_ctrl_5_s1_address                        => mm_interconnect_0_nco_freq_ctrl_5_s1_address,       --                          nco_freq_ctrl_5_s1.address
			nco_freq_ctrl_5_s1_write                          => mm_interconnect_0_nco_freq_ctrl_5_s1_write,         --                                            .write
			nco_freq_ctrl_5_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_5_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_5_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_5_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_5_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_5_s1_chipselect,    --                                            .chipselect
			nco_freq_ctrl_6_s1_address                        => mm_interconnect_0_nco_freq_ctrl_6_s1_address,       --                          nco_freq_ctrl_6_s1.address
			nco_freq_ctrl_6_s1_write                          => mm_interconnect_0_nco_freq_ctrl_6_s1_write,         --                                            .write
			nco_freq_ctrl_6_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_6_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_6_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_6_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_6_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_6_s1_chipselect,    --                                            .chipselect
			nco_freq_ctrl_7_s1_address                        => mm_interconnect_0_nco_freq_ctrl_7_s1_address,       --                          nco_freq_ctrl_7_s1.address
			nco_freq_ctrl_7_s1_write                          => mm_interconnect_0_nco_freq_ctrl_7_s1_write,         --                                            .write
			nco_freq_ctrl_7_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_7_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_7_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_7_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_7_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_7_s1_chipselect,    --                                            .chipselect
			nco_freq_ctrl_8_s1_address                        => mm_interconnect_0_nco_freq_ctrl_8_s1_address,       --                          nco_freq_ctrl_8_s1.address
			nco_freq_ctrl_8_s1_write                          => mm_interconnect_0_nco_freq_ctrl_8_s1_write,         --                                            .write
			nco_freq_ctrl_8_s1_readdata                       => mm_interconnect_0_nco_freq_ctrl_8_s1_readdata,      --                                            .readdata
			nco_freq_ctrl_8_s1_writedata                      => mm_interconnect_0_nco_freq_ctrl_8_s1_writedata,     --                                            .writedata
			nco_freq_ctrl_8_s1_chipselect                     => mm_interconnect_0_nco_freq_ctrl_8_s1_chipselect,    --                                            .chipselect
			nco_phase_ctrl_1_s1_address                       => mm_interconnect_0_nco_phase_ctrl_1_s1_address,      --                         nco_phase_ctrl_1_s1.address
			nco_phase_ctrl_1_s1_write                         => mm_interconnect_0_nco_phase_ctrl_1_s1_write,        --                                            .write
			nco_phase_ctrl_1_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_1_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_1_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_1_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_1_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_1_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_2_s1_address                       => mm_interconnect_0_nco_phase_ctrl_2_s1_address,      --                         nco_phase_ctrl_2_s1.address
			nco_phase_ctrl_2_s1_write                         => mm_interconnect_0_nco_phase_ctrl_2_s1_write,        --                                            .write
			nco_phase_ctrl_2_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_2_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_2_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_2_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_2_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_2_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_3_s1_address                       => mm_interconnect_0_nco_phase_ctrl_3_s1_address,      --                         nco_phase_ctrl_3_s1.address
			nco_phase_ctrl_3_s1_write                         => mm_interconnect_0_nco_phase_ctrl_3_s1_write,        --                                            .write
			nco_phase_ctrl_3_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_3_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_3_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_3_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_3_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_3_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_4_s1_address                       => mm_interconnect_0_nco_phase_ctrl_4_s1_address,      --                         nco_phase_ctrl_4_s1.address
			nco_phase_ctrl_4_s1_write                         => mm_interconnect_0_nco_phase_ctrl_4_s1_write,        --                                            .write
			nco_phase_ctrl_4_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_4_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_4_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_4_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_4_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_4_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_5_s1_address                       => mm_interconnect_0_nco_phase_ctrl_5_s1_address,      --                         nco_phase_ctrl_5_s1.address
			nco_phase_ctrl_5_s1_write                         => mm_interconnect_0_nco_phase_ctrl_5_s1_write,        --                                            .write
			nco_phase_ctrl_5_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_5_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_5_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_5_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_5_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_5_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_6_s1_address                       => mm_interconnect_0_nco_phase_ctrl_6_s1_address,      --                         nco_phase_ctrl_6_s1.address
			nco_phase_ctrl_6_s1_write                         => mm_interconnect_0_nco_phase_ctrl_6_s1_write,        --                                            .write
			nco_phase_ctrl_6_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_6_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_6_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_6_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_6_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_6_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_7_s1_address                       => mm_interconnect_0_nco_phase_ctrl_7_s1_address,      --                         nco_phase_ctrl_7_s1.address
			nco_phase_ctrl_7_s1_write                         => mm_interconnect_0_nco_phase_ctrl_7_s1_write,        --                                            .write
			nco_phase_ctrl_7_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_7_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_7_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_7_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_7_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_7_s1_chipselect,   --                                            .chipselect
			nco_phase_ctrl_8_s1_address                       => mm_interconnect_0_nco_phase_ctrl_8_s1_address,      --                         nco_phase_ctrl_8_s1.address
			nco_phase_ctrl_8_s1_write                         => mm_interconnect_0_nco_phase_ctrl_8_s1_write,        --                                            .write
			nco_phase_ctrl_8_s1_readdata                      => mm_interconnect_0_nco_phase_ctrl_8_s1_readdata,     --                                            .readdata
			nco_phase_ctrl_8_s1_writedata                     => mm_interconnect_0_nco_phase_ctrl_8_s1_writedata,    --                                            .writedata
			nco_phase_ctrl_8_s1_chipselect                    => mm_interconnect_0_nco_phase_ctrl_8_s1_chipselect,   --                                            .chipselect
			onchip_ram_s1_address                             => mm_interconnect_0_onchip_ram_s1_address,            --                               onchip_ram_s1.address
			onchip_ram_s1_write                               => mm_interconnect_0_onchip_ram_s1_write,              --                                            .write
			onchip_ram_s1_readdata                            => mm_interconnect_0_onchip_ram_s1_readdata,           --                                            .readdata
			onchip_ram_s1_writedata                           => mm_interconnect_0_onchip_ram_s1_writedata,          --                                            .writedata
			onchip_ram_s1_byteenable                          => mm_interconnect_0_onchip_ram_s1_byteenable,         --                                            .byteenable
			onchip_ram_s1_chipselect                          => mm_interconnect_0_onchip_ram_s1_chipselect,         --                                            .chipselect
			onchip_ram_s1_clken                               => mm_interconnect_0_onchip_ram_s1_clken               --                                            .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_nco_freq_control_1_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_control_1_s1_write;

	mm_interconnect_0_nco_freq_control_2_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_control_2_s1_write;

	mm_interconnect_0_nco_phase_ctrl_1_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_1_s1_write;

	mm_interconnect_0_nco_phase_ctrl_2_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_2_s1_write;

	mm_interconnect_0_gain_controller_s1_write_ports_inv <= not mm_interconnect_0_gain_controller_s1_write;

	mm_interconnect_0_nco_freq_ctrl_3_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_3_s1_write;

	mm_interconnect_0_nco_freq_ctrl_4_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_4_s1_write;

	mm_interconnect_0_nco_freq_ctrl_5_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_5_s1_write;

	mm_interconnect_0_nco_freq_ctrl_6_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_6_s1_write;

	mm_interconnect_0_nco_freq_ctrl_7_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_7_s1_write;

	mm_interconnect_0_nco_freq_ctrl_8_s1_write_ports_inv <= not mm_interconnect_0_nco_freq_ctrl_8_s1_write;

	mm_interconnect_0_nco_phase_ctrl_3_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_3_s1_write;

	mm_interconnect_0_nco_phase_ctrl_4_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_4_s1_write;

	mm_interconnect_0_nco_phase_ctrl_5_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_5_s1_write;

	mm_interconnect_0_nco_phase_ctrl_6_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_6_s1_write;

	mm_interconnect_0_nco_phase_ctrl_7_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_7_s1_write;

	mm_interconnect_0_nco_phase_ctrl_8_s1_write_ports_inv <= not mm_interconnect_0_nco_phase_ctrl_8_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of qsys_system
